package tdpram_tb_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;
	
	`include "tdpram_seq_item.svh"
	`include "tdpram_seq.svh"
	`include "tdpram_seqr.svh"
	`include "tdpram_drv.svh"
	`include "tdpram_cov.svh"
	`include "tdpram_mon1.svh"
	`include "tdpram_mon2.svh"
	`include "tdpram_agent1.svh"
	`include "tdpram_agent2.svh"
	`include "tdpram_sb.svh"
	`include "tdpram_env.svh"
	`include "tdpram_test.svh"
endpackage